** sch_path: /home/mona121130125/percobaan_layout/inverter_tb.sch
**.subckt inverter_tb
V1 net1 GND 1.8
V2 in GND PULSE(0 1.8 2NS 2NS 2NS 50NS 100NS 5)
x1 net1 in out GND inverter
**** begin user architecture code


.option wnflag=0
.option savecurrents
.control
save all
trans 1ns 200ns
plot in out
op
.endc


 .lib /home/mona121130125/pdk/sky130A/libs.tech/ngspice/models/sky130.lib.spice tt
.param mc_mm_switch=0
.param mc_pr_switch=1

**** end user architecture code
**.ends

* expanding   symbol:  /home/mona121130125/percobaan_layout/inverter.sym # of pins=4
** sym_path: /home/mona121130125/percobaan_layout/inverter.sym
** sch_path: /home/mona121130125/percobaan_layout/inverter.sch
.subckt inverter vdd in out gnd
*.ipin in
*.opin out
*.iopin vdd
*.iopin gnd
XM1 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
